`ifndef _TEST_TRANS_SVH
`define _TEST_TRANS_SVH

class test_transaction;
  bit [7:0] in;
  bit [7:0] out;
endclass

`endif
